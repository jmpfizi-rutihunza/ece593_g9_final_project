package mp_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "mp_seq_item.sv"
  `include "mp_driver.sv"
  `include "mp_req_monitor.sv"
  `include "mp_rsp_monitor.sv"
  `include "mp_scoreboard.sv"
  `include "mp_agent.sv"
  `include "mp_env.sv"
  `include "mp_test.sv"

endpackage
