//////////////////////////////////////////////////
//  ECE-593 Project                              //
//  Multiprocessor System                        //
//  Milestone2 - Functional Coverage             //
//////////////////////////////////////////////////

`include "transaction.sv"

class coverage;

  // Covergroup sampled via function call (tool-friendly & simple)
  covergroup cg_tr with function sample(
      bit [1:0]  core_id,
      bit [3:0]  opcode,
      bit [10:0] addr,
      bit        we
  );

    // Which core issued the transaction
    cp_core: coverpoint core_id {
      bins c0 = {2'd0};
      bins c1 = {2'd1};
      bins c2 = {2'd2};
      bins c3 = {2'd3};
    }

    // Opcode coverage (bins for your valid range)
    cp_opcode: coverpoint opcode {
      bins op_valid[] = {[4'h0:4'hD]};
      illegal_bins op_illegal = default;
    }

    // Address space partitioning (2KB memory => addr < 2048)
    cp_addr: coverpoint addr {
      bins low  = {[11'd0   : 11'd255]};
      bins mid  = {[11'd256 : 11'd1023]};
      bins high = {[11'd1024: 11'd2047]};
      illegal_bins bad = default;
    }

    // Read vs write (based on we)
    cp_we: coverpoint we {
      bins read  = {1'b0};
      bins write = {1'b1};
    }

    // Crosses (these are usually what graders like seeing)
    x_core_opcode : cross cp_core, cp_opcode;
    x_we_opcode   : cross cp_we,   cp_opcode;

  endgroup

  function new();
    cg_tr = new();
  endfunction

  // call this from SCB (or monitor) on real observed transactions
  function void sample(transaction t);
    cg_tr.sample(t.core_id, t.opcode, t.addr, t.we);
  endfunction

endclass
