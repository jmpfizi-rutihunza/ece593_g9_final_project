package tb_pkg;

   `include "transaction.sv"
   `include "coverage_collector.sv"

endpackage